module direction();
 
endmodule 